`ifndef module_SD
`define module_SD

`include "config/config.sv"

module SD(

);

endmodule

`endif
