`timescale 1ns/1ps

`include "lab08.sv"

module RAM_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

RAM tb(

);

endmodule

