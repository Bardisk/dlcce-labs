`timescale 1ns/1ps

`include "lab11.sv"

module lab11_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

lab11 tb(

);

endmodule

