`ifndef module_Memory
`define module_Memory

`include "config/config.sv"

module Memory(

);

endmodule

`endif
