`timescale 1ns/1ps

`include "lab07.sv"

module debounce_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

debounce tb(

);

endmodule

