`timescale 1ns/1ps

`include "lab11.sv"

module inst_memory_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

inst_memory tb(

);

endmodule

