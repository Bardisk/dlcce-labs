`ifndef module_template
`define module_template

`include "config/config.sv"

module template(

);

endmodule

`endif
