`define SIM

`include "config/config.sv"
//add includes here

module template(
 
);


endmodule
