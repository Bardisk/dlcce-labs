`ifndef module_debounce
`define module_debounce

module debounce(
    
);

endmodule

`endif
