`ifndef module_ledTubes
`define module_ledTubes

`include "ledTubes/ledTube.sv"
`include "ledTubes/timeoutledTube.sv"

`endif
