module template(

);

endmodule