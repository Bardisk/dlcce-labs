`define SIM

`include "ledmonitor/ledmonitor.sv"
`include "clockGenerator/clockGenerator.sv"
`include "regfile/regfile.sv"
//add includes here

module lab05(
 
);


endmodule
