`timescale 1ns/1ps

`include "unisys.sv"

module VGA_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

VGA tb(

);

endmodule

