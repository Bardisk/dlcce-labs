`timescale 1ns/1ps

`include "unisys.sv"

module Memory_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

Memory tb(

);

endmodule

