`timescale 1ns/1ps

`include "lab11.sv"

module Bus_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

Bus tb(

);

endmodule

