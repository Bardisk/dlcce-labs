`ifndef module_VGA
`define module_VGA

`include "config/config.sv"

module VGA(

);

endmodule

`endif
