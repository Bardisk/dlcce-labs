`timescale 1ns/1ps

`include "lab11.sv"

module ALU_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

ALU tb(

);

endmodule

