`timescale 1ns/1ps

`include "lab07.sv"

module keyboardCtr_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

keyboardCtr tb(

);

endmodule

