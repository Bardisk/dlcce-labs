`define SIM

`include "clockGenerator/clockGenerator.sv"
`include "RAM/RAM.sv"
`include "Visual_Adapter/Visual_Adapter.sv"
`include "keyboardCtr/keyboardCtr.sv"
`include "Simple_Bus/Simple_Bus.sv"
`include "Vga_Ctr/Vga_Ctr.sv"
`include "ledmonitor/ledmonitor.sv"
`include "config/config.sv"
//add includes here

module lab09(
 
);


endmodule
