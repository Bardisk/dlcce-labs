`ifndef module_CPU
`define module_CPU

`include "config/config.sv"

module CPU(

);

endmodule

`endif
