`timescale 1ns/1ps

`include "lab07.sv"

module lab07_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

lab07 tb(

);

endmodule

