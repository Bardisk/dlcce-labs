`define SIM

//add includes here

module template(
 
);


endmodule
