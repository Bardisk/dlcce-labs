`ifndef module_Timer
`define module_Timer

`include "config/config.sv"

module Timer(

);

endmodule

`endif
