`timescale 1ns/1ps

`include "lab09.sv"

module lab09_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

lab09 tb(

);

endmodule

