`ifndef module_Keyboard
`define module_Keyboard

`include "config/config.sv"

module Keyboard(

);

endmodule

`endif
