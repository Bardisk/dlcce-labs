`define SIM

`include "config/config.sv"
`include "control_signal_generator/control_signal_generator.sv"
`include "imm_generator/imm_generator.sv"
`include "pc_generator/pc_generator.sv"
`include "inst_memory/inst_memory.sv"
`include "data_memory/data_memory.sv"
`include "regheap/regheap.sv"
`include "CPU/CPU.sv"
`include "ALU/ALU.sv"
`include "jump_control/jump_control.sv"
`include "Bus/Bus.sv"
`include "ojcpu/ojcpu.sv"
//add includes here

module lab11(
 
);


endmodule
