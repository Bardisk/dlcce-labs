`timescale 1ns/1ps

`include "lab09.sv"

module Kbd_CU_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

Kbd_CU tb(

);

endmodule

