`timescale 1ns/1ps

`include "lab05.sv"

module regfile_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

regfile tb(

);

endmodule

