`ifndef module_Number_Screen
`define module_Number_Screen

`include "config/config.sv"

module Number_Screen(

);

endmodule

`endif
