`timescale 1ns/1ps

`include "lab07.sv"

module codeToAscii_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

codeToAscii tb(

);

endmodule

