`timescale 1ns/1ps

`include "unisys.sv"

module Keyboard_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

Keyboard tb(

);

endmodule

