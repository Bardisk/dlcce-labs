`timescale 1ns/1ps

`include "unisys.sv"

module SIB_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

SIB tb(

);

endmodule

