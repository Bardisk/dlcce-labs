`timescale 1ns/1ps

`include "unisys.sv"

module Timer_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

Timer tb(

);

endmodule

