`timescale 1ns/1ps

`include "lab11.sv"

module imm_generator_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

imm_generator tb(

);

endmodule

