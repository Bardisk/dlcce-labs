`ifndef module_Simple_Bus
`define module_Simple_Bus

module Simple_Bus(

);

endmodule

`endif
