`ifndef module_template
`define module_template

module template(

);

endmodule

`endif
