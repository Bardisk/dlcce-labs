`ifndef module_memory_config
`define module_memory_config

`define MAIN_ADDR_WIDTH 18
`define MAIN_ADDR_WIDE  `MAIN_ADDR_WIDTH:0
`define VGM_ADDR_WIDTH  18
`define VCM_ADDR_WIDTH  13
`define VGM_SIZE        307200
`define VCM_SIZE        2100
`define VGM_WIDTH       4
`define VCM_WIDTH       12
`define VGM_WIDE        `VGM_WIDTH-1:0
`define VCM_WIDE        `VCM_WIDTH-1:0

`VGA_

`endif
