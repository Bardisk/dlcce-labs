`ifndef module_SIB
`define module_SIB

`include "config/config.sv"

module SIB(

);

endmodule

`endif
