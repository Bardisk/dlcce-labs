`timescale 1ns/1ps

`include "lab11.sv"

module control_signal_generator_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

control_signal_generator tb(

);

endmodule

