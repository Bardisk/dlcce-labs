`timescale 1ns/1ps

`include "encryption.sv"

module encryption_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

encryption tb(

);

endmodule

