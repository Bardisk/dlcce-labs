`timescale 1ns/1ps

`include "unisys.sv"

module CPU_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

CPU tb(

);

endmodule

