`timescale 1ns/1ps

`include "lab07.sv"

module ps2Keyboard_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

ps2Keyboard tb(

);

endmodule

