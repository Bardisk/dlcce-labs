`timescale 1ns/1ps

`include "lab11.sv"

module regheap_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

regheap tb(

);

endmodule

