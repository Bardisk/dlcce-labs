`timescale 1ns/1ps

`include "lab08.sv"

module Mem_Ctr_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

Mem_Ctr tb(

);

endmodule

