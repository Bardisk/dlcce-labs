`timescale 1ns/1ps

`include "lab11.sv"

module data_memory_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

data_memory tb(

);

endmodule

