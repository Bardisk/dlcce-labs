module template(

);

endmodule
