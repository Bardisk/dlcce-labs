`timescale 1ns/1ps

`include "lab05.sv"

module lab05_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

lab05 tb(

);

endmodule

