`timescale 1ns/1ps

`include "lab11.sv"

module jump_control_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

jump_control tb(

);

endmodule

