`timescale 1ns/1ps

`include "unisys.sv"

module SD_tb();

initial begin
    $dumpfile("build/wave.vcd");
    $dumpvars;
end

SD tb(

);

endmodule

